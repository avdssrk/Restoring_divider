`timescale 1ns / 1ps

module test_bench();
    //test bench for divider
    reg [7:0] n,d;
    
    wire [7:0] q;
    Divd uut(n,d,q);
    initial begin
        n=8'b1000_0000;  //8
        d=8'b1111_0000;  //15
        
        #100
        n=8'b0100_0000;  //8
        d=8'b0000_1000;  //0.5
        
        #100
        n=8'b1010_0000;  //10
        d=8'b0101_0000;  //5
        
        #100
        n=8'b1000_1000;  //8.5
        d=8'b0010_0000;  //2
        
        #100
        n=8'b0010_0000;  //2
        d=8'b0011_0000;  //3
        
        #100
        n=8'b0010_0000;  //2
        d=8'b0100_0000;  //4
        
        #100 
        n = 8'b0001_0000; //1
        d = 8'b0010_0000; //2
        
        
    end
       
    
endmodule
